module q1_3(a,f);
input a;
output f;
assign f = ~(~a);
endmodule
